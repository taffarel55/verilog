module hello;
initial
begin
    $display("Hello word!");
    $finish;
end
endmodule