module or2(
    output y,
    input a,b
);

assign y = a | b;

endmodule